`timescale 1ns / 1ps

module decoder(in_char1, in_char2, char1, char2);
	input [3:0] in_char1, in_char2; 
	output [3:0] char1, char2; 

	reg [3:0] char1, char1;
	
	assign char1 = char1 - 1;
    assign char2 = char2 - 1;
endmodule